library verilog;
use verilog.vl_types.all;
entity ConditionalLogic_vlg_vec_tst is
end ConditionalLogic_vlg_vec_tst;
