library verilog;
use verilog.vl_types.all;
entity topmodule_vlg_vec_tst is
end topmodule_vlg_vec_tst;
